-- Superawesome Project Processor

entity toplevel is
	-- Generics
	-- Ports
end entity;

architecture behaviour of toplevel is
	-- Components
begin
	-- Instantiations
end behaviour;


entity core is
	-- Generics
	-- Ports
end entity;

architecture behaviour of core is
	-- Components
begin
	-- Instantiations
end behaviour;

entity EBI is
	-- Generics
	-- Ports
end entity;

architecture behaviour of EBI is
	-- Components
begin
	-- Instantiations
end behaviour;

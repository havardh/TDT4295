entity pipeline is
	-- Generics
	-- Ports
end entity;

architecture behaviour of pipeline is
	-- Components
begin
	-- Instantiations
end behaviour;

entity procbuffer is
	-- Generics
	-- Ports
end entity;

architecture behaviour of procbuffer is
	-- Components
begin
	-- Instantiations
end behaviour;

entity processorcore is
	-- Generics
	-- Ports
end entity;

architecture behaviour of processorcore is
	-- Components
begin
	-- Instantiations
end behaviour;
